-- Trabajo SED 23/24 Grupo 2
-- Modulo display
-- Entidad de configuración de la
-- visualizacion en formato 12h/24h


--entity display is
--    Port (
--        CLK100MHZ  : in std_logic;
--        mode: in std_logic_vector(3 downto 0);
--        buttons: in std_logic_vector(3 downto 0);
--        digits_0to3 : in std_logic_vector(15 downto 0);
--        digits_4to7 : in std_logic_vector(15 downto 0);
--        blink_pairs : in std_logic_vector(3 downto 0);
--        out_mode : out std_logic_vector(3 downto 0)
--    );
--end display;




--architecture Behavioral of display is
--begin
--	out_mode <= '1' when (buttons = "1000" and mode = "1000") else unaffected;
--	out_mode <= '0' when (buttons = "0010" and mode = "1000") else unaffected;
	
--	digits_0to3 <= 
--end Behavioral;


